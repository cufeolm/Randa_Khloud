`include "add.svh"
`include "test.svh"
`include "swap.svh"
`include "swap_byte.svh"
`include "swap_ans.svh"
`include "set_high_order.svh"
`include "atomic_load_store.svh"
`include "atomic_load_store_ans.svh"
`include "load_s_byte.svh"
`include "load_u_byte.svh"